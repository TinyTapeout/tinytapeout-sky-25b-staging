module tt_um_technology_characterization (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire chain_out;
 wire \clkgen_inst.cnt_1m[0] ;
 wire \clkgen_inst.cnt_1m[1] ;
 wire \clkgen_inst.cnt_1m[2] ;
 wire \clkgen_inst.cnt_1m[3] ;
 wire \clkgen_inst.cnt_1m[4] ;
 wire \clkgen_inst.cnt_1m[5] ;
 wire \clkgen_inst.cnt_1s[0] ;
 wire \clkgen_inst.cnt_1s[10] ;
 wire \clkgen_inst.cnt_1s[11] ;
 wire \clkgen_inst.cnt_1s[12] ;
 wire \clkgen_inst.cnt_1s[13] ;
 wire \clkgen_inst.cnt_1s[14] ;
 wire \clkgen_inst.cnt_1s[15] ;
 wire \clkgen_inst.cnt_1s[16] ;
 wire \clkgen_inst.cnt_1s[17] ;
 wire \clkgen_inst.cnt_1s[18] ;
 wire \clkgen_inst.cnt_1s[19] ;
 wire \clkgen_inst.cnt_1s[1] ;
 wire \clkgen_inst.cnt_1s[20] ;
 wire \clkgen_inst.cnt_1s[21] ;
 wire \clkgen_inst.cnt_1s[22] ;
 wire \clkgen_inst.cnt_1s[23] ;
 wire \clkgen_inst.cnt_1s[24] ;
 wire \clkgen_inst.cnt_1s[25] ;
 wire \clkgen_inst.cnt_1s[2] ;
 wire \clkgen_inst.cnt_1s[3] ;
 wire \clkgen_inst.cnt_1s[4] ;
 wire \clkgen_inst.cnt_1s[5] ;
 wire \clkgen_inst.cnt_1s[6] ;
 wire \clkgen_inst.cnt_1s[7] ;
 wire \clkgen_inst.cnt_1s[8] ;
 wire \clkgen_inst.cnt_1s[9] ;
 wire \clkgen_inst.htol_1Mhz_toggle ;
 wire \clkgen_inst.htol_1s_toggle ;
 wire \clkgen_inst.n28_o[0] ;
 wire \clkgen_inst.n28_o[10] ;
 wire \clkgen_inst.n28_o[11] ;
 wire \clkgen_inst.n28_o[12] ;
 wire \clkgen_inst.n28_o[13] ;
 wire \clkgen_inst.n28_o[14] ;
 wire \clkgen_inst.n28_o[15] ;
 wire \clkgen_inst.n28_o[16] ;
 wire \clkgen_inst.n28_o[17] ;
 wire \clkgen_inst.n28_o[18] ;
 wire \clkgen_inst.n28_o[19] ;
 wire \clkgen_inst.n28_o[1] ;
 wire \clkgen_inst.n28_o[20] ;
 wire \clkgen_inst.n28_o[21] ;
 wire \clkgen_inst.n28_o[22] ;
 wire \clkgen_inst.n28_o[23] ;
 wire \clkgen_inst.n28_o[24] ;
 wire \clkgen_inst.n28_o[25] ;
 wire \clkgen_inst.n28_o[2] ;
 wire \clkgen_inst.n28_o[3] ;
 wire \clkgen_inst.n28_o[4] ;
 wire \clkgen_inst.n28_o[5] ;
 wire \clkgen_inst.n28_o[6] ;
 wire \clkgen_inst.n28_o[7] ;
 wire \clkgen_inst.n28_o[8] ;
 wire \clkgen_inst.n28_o[9] ;
 wire \clkgen_inst.n30_o[0] ;
 wire \clkgen_inst.n30_o[1] ;
 wire \clkgen_inst.n30_o[2] ;
 wire \clkgen_inst.n30_o[3] ;
 wire \clkgen_inst.n30_o[4] ;
 wire \clkgen_inst.n30_o[5] ;
 wire htol_latched;
 wire \inverterchain_inst.chain_3q ;
 wire \inverterchain_inst.chain_mid ;
 wire \inverterchain_inst.gen_inv_n1000_inv_inst.A ;
 wire \inverterchain_inst.gen_inv_n1000_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1001_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1002_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1003_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1004_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1005_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1006_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1007_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1008_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1009_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n100_inv_inst.A ;
 wire \inverterchain_inst.gen_inv_n100_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1010_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1011_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1012_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1013_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1014_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1015_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1016_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1017_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1018_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1019_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n101_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1020_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1021_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1022_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1023_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n102_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n103_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n104_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n105_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n106_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n107_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n108_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n109_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n10_inv_inst.A ;
 wire \inverterchain_inst.gen_inv_n10_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n110_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n111_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n112_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n113_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n114_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n115_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n116_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n117_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n118_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n119_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n11_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n120_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n121_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n122_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n123_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n124_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n125_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n126_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n127_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n128_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n129_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n12_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n130_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n131_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n132_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n133_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n134_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n135_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n136_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n137_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n138_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n139_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n13_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n140_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n141_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n142_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n143_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n144_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n145_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n146_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n147_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n148_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n149_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n14_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n150_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n151_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n152_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n153_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n154_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n155_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n156_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n157_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n158_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n159_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n15_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n160_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n161_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n162_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n163_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n164_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n165_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n166_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n167_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n168_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n169_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n16_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n170_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n171_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n172_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n173_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n174_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n175_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n176_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n177_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n178_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n179_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n17_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n180_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n181_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n182_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n183_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n184_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n185_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n186_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n187_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n188_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n189_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n18_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n190_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n191_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n192_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n193_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n194_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n195_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n196_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n197_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n198_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n199_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n19_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n1_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n200_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n201_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n202_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n203_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n204_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n205_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n206_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n207_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n208_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n209_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n20_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n210_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n211_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n212_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n213_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n214_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n215_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n216_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n217_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n218_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n219_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n21_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n220_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n221_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n222_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n223_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n224_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n225_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n226_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n227_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n228_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n229_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n22_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n230_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n231_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n232_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n233_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n234_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n235_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n236_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n237_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n238_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n239_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n23_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n240_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n241_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n242_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n243_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n244_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n245_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n246_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n247_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n248_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n249_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n24_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n250_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n251_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n252_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n253_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n254_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n255_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n256_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n257_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n258_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n259_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n25_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n260_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n261_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n262_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n263_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n264_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n265_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n266_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n267_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n268_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n269_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n26_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n270_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n271_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n272_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n273_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n274_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n275_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n276_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n277_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n278_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n279_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n27_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n280_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n281_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n282_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n283_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n284_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n285_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n286_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n287_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n288_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n289_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n28_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n290_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n291_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n292_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n293_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n294_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n295_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n296_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n297_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n298_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n299_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n29_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n2_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n300_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n301_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n302_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n303_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n304_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n305_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n306_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n307_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n308_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n309_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n30_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n310_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n311_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n312_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n313_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n314_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n315_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n316_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n317_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n318_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n319_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n31_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n320_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n321_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n322_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n323_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n324_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n325_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n326_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n327_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n328_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n329_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n32_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n330_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n331_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n332_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n333_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n334_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n335_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n336_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n337_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n338_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n339_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n33_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n340_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n341_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n342_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n343_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n344_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n345_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n346_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n347_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n348_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n349_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n34_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n350_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n351_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n352_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n353_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n354_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n355_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n356_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n357_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n358_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n359_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n35_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n360_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n361_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n362_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n363_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n364_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n365_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n366_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n367_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n368_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n369_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n36_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n370_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n371_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n372_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n373_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n374_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n375_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n376_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n377_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n378_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n379_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n37_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n380_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n381_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n382_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n383_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n384_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n385_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n386_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n387_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n388_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n389_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n38_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n390_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n391_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n392_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n393_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n394_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n395_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n396_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n397_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n398_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n399_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n39_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n3_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n400_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n401_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n402_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n403_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n404_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n405_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n406_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n407_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n408_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n409_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n40_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n410_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n411_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n412_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n413_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n414_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n415_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n416_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n417_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n418_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n419_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n41_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n420_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n421_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n422_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n423_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n424_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n425_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n426_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n427_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n428_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n429_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n42_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n430_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n431_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n432_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n433_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n434_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n435_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n436_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n437_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n438_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n439_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n43_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n440_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n441_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n442_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n443_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n444_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n445_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n446_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n447_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n448_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n449_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n44_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n450_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n451_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n452_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n453_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n454_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n455_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n456_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n457_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n458_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n459_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n45_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n460_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n461_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n462_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n463_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n464_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n465_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n466_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n467_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n468_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n469_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n46_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n470_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n471_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n472_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n473_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n474_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n475_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n476_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n477_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n478_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n479_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n47_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n480_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n481_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n482_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n483_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n484_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n485_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n486_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n487_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n488_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n489_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n48_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n490_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n491_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n492_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n493_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n494_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n495_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n496_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n497_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n498_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n499_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n49_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n4_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n500_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n501_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n502_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n503_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n504_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n505_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n506_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n507_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n508_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n509_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n50_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n510_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n511_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n513_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n514_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n515_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n516_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n517_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n518_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n519_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n51_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n520_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n521_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n522_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n523_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n524_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n525_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n526_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n527_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n528_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n529_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n52_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n530_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n531_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n532_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n533_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n534_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n535_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n536_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n537_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n538_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n539_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n53_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n540_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n541_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n542_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n543_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n544_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n545_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n546_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n547_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n548_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n549_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n54_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n550_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n551_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n552_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n553_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n554_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n555_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n556_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n557_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n558_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n559_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n55_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n560_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n561_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n562_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n563_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n564_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n565_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n566_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n567_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n568_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n569_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n56_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n570_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n571_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n572_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n573_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n574_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n575_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n576_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n577_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n578_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n579_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n57_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n580_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n581_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n582_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n583_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n584_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n585_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n586_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n587_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n588_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n589_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n58_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n590_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n591_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n592_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n593_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n594_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n595_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n596_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n597_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n598_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n599_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n59_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n5_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n600_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n601_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n602_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n603_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n604_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n605_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n606_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n607_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n608_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n609_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n60_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n610_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n611_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n612_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n613_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n614_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n615_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n616_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n617_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n618_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n619_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n61_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n620_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n621_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n622_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n623_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n624_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n625_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n626_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n627_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n628_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n629_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n62_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n630_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n631_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n632_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n633_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n634_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n635_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n636_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n637_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n638_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n639_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n63_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n640_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n641_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n642_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n643_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n644_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n645_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n646_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n647_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n648_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n649_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n64_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n650_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n651_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n652_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n653_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n654_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n655_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n656_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n657_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n658_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n659_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n65_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n660_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n661_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n662_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n663_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n664_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n665_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n666_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n667_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n668_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n669_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n66_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n670_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n671_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n672_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n673_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n674_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n675_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n676_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n677_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n678_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n679_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n67_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n680_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n681_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n682_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n683_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n684_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n685_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n686_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n687_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n688_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n689_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n68_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n690_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n691_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n692_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n693_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n694_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n695_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n696_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n697_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n698_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n699_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n69_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n6_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n700_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n701_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n702_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n703_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n704_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n705_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n706_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n707_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n708_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n709_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n70_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n710_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n711_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n712_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n713_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n714_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n715_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n716_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n717_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n718_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n719_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n71_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n720_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n721_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n722_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n723_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n724_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n725_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n726_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n727_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n728_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n729_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n72_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n730_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n731_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n732_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n733_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n734_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n735_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n736_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n737_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n738_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n739_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n73_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n740_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n741_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n742_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n743_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n744_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n745_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n746_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n747_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n748_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n749_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n74_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n750_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n751_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n752_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n753_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n754_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n755_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n756_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n757_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n758_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n759_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n75_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n760_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n761_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n762_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n763_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n764_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n765_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n766_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n767_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n769_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n76_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n770_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n771_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n772_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n773_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n774_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n775_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n776_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n777_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n778_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n779_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n77_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n780_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n781_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n782_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n783_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n784_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n785_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n786_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n787_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n788_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n789_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n78_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n790_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n791_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n792_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n793_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n794_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n795_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n796_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n797_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n798_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n799_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n79_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n7_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n800_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n801_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n802_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n803_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n804_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n805_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n806_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n807_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n808_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n809_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n80_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n810_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n811_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n812_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n813_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n814_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n815_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n816_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n817_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n818_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n819_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n81_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n820_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n821_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n822_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n823_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n824_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n825_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n826_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n827_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n828_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n829_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n82_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n830_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n831_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n832_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n833_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n834_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n835_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n836_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n837_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n838_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n839_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n83_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n840_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n841_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n842_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n843_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n844_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n845_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n846_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n847_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n848_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n849_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n84_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n850_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n851_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n852_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n853_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n854_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n855_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n856_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n857_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n858_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n859_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n85_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n860_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n861_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n862_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n863_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n864_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n865_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n866_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n867_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n868_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n869_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n86_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n870_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n871_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n872_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n873_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n874_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n875_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n876_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n877_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n878_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n879_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n87_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n880_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n881_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n882_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n883_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n884_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n885_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n886_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n887_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n888_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n889_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n88_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n890_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n891_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n892_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n893_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n894_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n895_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n896_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n897_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n898_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n899_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n89_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n8_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n900_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n901_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n902_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n903_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n904_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n905_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n906_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n907_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n908_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n909_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n90_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n910_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n911_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n912_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n913_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n914_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n915_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n916_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n917_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n918_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n919_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n91_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n920_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n921_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n922_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n923_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n924_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n925_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n926_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n927_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n928_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n929_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n92_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n930_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n931_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n932_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n933_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n934_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n935_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n936_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n937_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n938_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n939_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n93_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n940_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n941_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n942_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n943_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n944_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n945_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n946_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n947_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n948_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n949_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n94_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n950_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n951_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n952_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n953_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n954_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n955_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n956_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n957_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n958_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n959_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n95_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n960_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n961_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n962_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n963_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n964_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n965_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n966_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n967_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n968_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n969_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n96_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n970_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n971_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n972_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n973_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n974_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n975_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n976_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n977_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n978_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n979_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n97_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n980_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n981_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n982_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n983_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n984_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n985_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n986_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n987_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n988_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n989_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n98_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n990_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n991_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n992_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n993_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n994_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n995_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n996_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n997_inv_inst.Y ;
 wire \inverterchain_inst.gen_inv_n998_inv_inst.Y ;
 wire n55_o;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;

 sky130_fd_sc_hd__inv_2 _082_ (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _083_ (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _084_ (.A(\clkgen_inst.cnt_1s[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _085_ (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _086_ (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _087_ (.A(net9),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _088_ (.A(\clkgen_inst.htol_1Mhz_toggle ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_077_));
 sky130_fd_sc_hd__or3_1 _089_ (.A(net7),
    .B(net6),
    .C(htol_latched),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_078_));
 sky130_fd_sc_hd__a2111oi_4 _090_ (.A1(net5),
    .A2(_076_),
    .B1(_078_),
    .C1(net4),
    .D1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(uo_out[4]));
 sky130_fd_sc_hd__a21o_2 _091_ (.A1(net17),
    .A2(htol_latched),
    .B1(uo_out[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[5]));
 sky130_fd_sc_hd__a31o_4 _092_ (.A1(net17),
    .A2(htol_latched),
    .A3(\clkgen_inst.htol_1Mhz_toggle ),
    .B1(uo_out[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[6]));
 sky130_fd_sc_hd__a31o_2 _093_ (.A1(net17),
    .A2(htol_latched),
    .A3(clknet_2_1__leaf_clk),
    .B1(uo_out[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[7]));
 sky130_fd_sc_hd__nand2b_1 _094_ (.A_N(\clkgen_inst.htol_1s_toggle ),
    .B(htol_latched),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n55_o));
 sky130_fd_sc_hd__or2_1 _095_ (.A(\clkgen_inst.cnt_1m[1] ),
    .B(\clkgen_inst.cnt_1m[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_079_));
 sky130_fd_sc_hd__nand2_1 _096_ (.A(\clkgen_inst.cnt_1m[3] ),
    .B(\clkgen_inst.cnt_1m[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_080_));
 sky130_fd_sc_hd__or4_1 _097_ (.A(\clkgen_inst.cnt_1m[2] ),
    .B(\clkgen_inst.cnt_1m[5] ),
    .C(_079_),
    .D(_080_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_081_));
 sky130_fd_sc_hd__and2_1 _098_ (.A(net17),
    .B(_081_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_003_));
 sky130_fd_sc_hd__and2b_1 _099_ (.A_N(\clkgen_inst.cnt_1m[0] ),
    .B(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n30_o[0] ));
 sky130_fd_sc_hd__nand2_1 _100_ (.A(\clkgen_inst.cnt_1m[1] ),
    .B(\clkgen_inst.cnt_1m[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_004_));
 sky130_fd_sc_hd__and3_1 _101_ (.A(net17),
    .B(_079_),
    .C(_004_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n30_o[1] ));
 sky130_fd_sc_hd__a21o_1 _102_ (.A1(\clkgen_inst.cnt_1m[1] ),
    .A2(\clkgen_inst.cnt_1m[0] ),
    .B1(\clkgen_inst.cnt_1m[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_005_));
 sky130_fd_sc_hd__and3_1 _103_ (.A(\clkgen_inst.cnt_1m[1] ),
    .B(\clkgen_inst.cnt_1m[0] ),
    .C(\clkgen_inst.cnt_1m[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_006_));
 sky130_fd_sc_hd__and3b_1 _104_ (.A_N(_006_),
    .B(net17),
    .C(_005_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n30_o[2] ));
 sky130_fd_sc_hd__and2_1 _105_ (.A(\clkgen_inst.cnt_1m[3] ),
    .B(_006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_007_));
 sky130_fd_sc_hd__o21ai_1 _106_ (.A1(net48),
    .A2(_006_),
    .B1(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_008_));
 sky130_fd_sc_hd__nor2_1 _107_ (.A(_007_),
    .B(_008_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n30_o[3] ));
 sky130_fd_sc_hd__and3_1 _108_ (.A(\clkgen_inst.cnt_1m[3] ),
    .B(\clkgen_inst.cnt_1m[4] ),
    .C(_006_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_009_));
 sky130_fd_sc_hd__inv_2 _109_ (.A(_009_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_010_));
 sky130_fd_sc_hd__o211a_1 _110_ (.A1(net41),
    .A2(_007_),
    .B1(_010_),
    .C1(_003_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n30_o[4] ));
 sky130_fd_sc_hd__o21ai_1 _111_ (.A1(net37),
    .A2(_009_),
    .B1(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_011_));
 sky130_fd_sc_hd__a21oi_1 _112_ (.A1(net37),
    .A2(_009_),
    .B1(_011_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n30_o[5] ));
 sky130_fd_sc_hd__nor2_1 _113_ (.A(net12),
    .B(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n28_o[0] ));
 sky130_fd_sc_hd__a21oi_1 _114_ (.A1(\clkgen_inst.cnt_1s[1] ),
    .A2(\clkgen_inst.cnt_1s[0] ),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_012_));
 sky130_fd_sc_hd__o21a_1 _115_ (.A1(\clkgen_inst.cnt_1s[1] ),
    .A2(net38),
    .B1(_012_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[1] ));
 sky130_fd_sc_hd__a21oi_1 _116_ (.A1(\clkgen_inst.cnt_1s[1] ),
    .A2(\clkgen_inst.cnt_1s[0] ),
    .B1(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_013_));
 sky130_fd_sc_hd__a31o_1 _117_ (.A1(\clkgen_inst.cnt_1s[1] ),
    .A2(\clkgen_inst.cnt_1s[0] ),
    .A3(\clkgen_inst.cnt_1s[2] ),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_014_));
 sky130_fd_sc_hd__nor2_1 _118_ (.A(_013_),
    .B(_014_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n28_o[2] ));
 sky130_fd_sc_hd__a31o_1 _119_ (.A1(\clkgen_inst.cnt_1s[1] ),
    .A2(\clkgen_inst.cnt_1s[0] ),
    .A3(\clkgen_inst.cnt_1s[2] ),
    .B1(\clkgen_inst.cnt_1s[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_015_));
 sky130_fd_sc_hd__and4_2 _120_ (.A(\clkgen_inst.cnt_1s[1] ),
    .B(\clkgen_inst.cnt_1s[0] ),
    .C(\clkgen_inst.cnt_1s[3] ),
    .D(\clkgen_inst.cnt_1s[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_016_));
 sky130_fd_sc_hd__and3b_1 _121_ (.A_N(_016_),
    .B(net18),
    .C(_015_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[3] ));
 sky130_fd_sc_hd__a21oi_1 _122_ (.A1(\clkgen_inst.cnt_1s[4] ),
    .A2(_016_),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_017_));
 sky130_fd_sc_hd__o21a_1 _123_ (.A1(\clkgen_inst.cnt_1s[4] ),
    .A2(_016_),
    .B1(_017_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[4] ));
 sky130_fd_sc_hd__a21o_1 _124_ (.A1(\clkgen_inst.cnt_1s[4] ),
    .A2(_016_),
    .B1(\clkgen_inst.cnt_1s[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_018_));
 sky130_fd_sc_hd__and3_1 _125_ (.A(\clkgen_inst.cnt_1s[5] ),
    .B(\clkgen_inst.cnt_1s[4] ),
    .C(_016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_019_));
 sky130_fd_sc_hd__nand3_1 _126_ (.A(\clkgen_inst.cnt_1s[5] ),
    .B(\clkgen_inst.cnt_1s[4] ),
    .C(_016_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_020_));
 sky130_fd_sc_hd__and3_1 _127_ (.A(net17),
    .B(_018_),
    .C(_020_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[5] ));
 sky130_fd_sc_hd__or4bb_1 _128_ (.A(\clkgen_inst.cnt_1s[23] ),
    .B(\clkgen_inst.cnt_1s[25] ),
    .C_N(\clkgen_inst.cnt_1s[24] ),
    .D_N(\clkgen_inst.cnt_1s[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_021_));
 sky130_fd_sc_hd__nand2_1 _129_ (.A(\clkgen_inst.cnt_1s[14] ),
    .B(\clkgen_inst.cnt_1s[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_022_));
 sky130_fd_sc_hd__or4b_1 _130_ (.A(\clkgen_inst.cnt_1s[9] ),
    .B(\clkgen_inst.cnt_1s[8] ),
    .C(\clkgen_inst.cnt_1s[10] ),
    .D_N(\clkgen_inst.cnt_1s[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_023_));
 sky130_fd_sc_hd__or4_1 _131_ (.A(\clkgen_inst.cnt_1s[15] ),
    .B(\clkgen_inst.cnt_1s[17] ),
    .C(_022_),
    .D(_023_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_024_));
 sky130_fd_sc_hd__and2_1 _132_ (.A(\clkgen_inst.cnt_1s[13] ),
    .B(\clkgen_inst.cnt_1s[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_025_));
 sky130_fd_sc_hd__and2_1 _133_ (.A(\clkgen_inst.cnt_1s[21] ),
    .B(\clkgen_inst.cnt_1s[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_026_));
 sky130_fd_sc_hd__nand4_1 _134_ (.A(\clkgen_inst.cnt_1s[13] ),
    .B(\clkgen_inst.cnt_1s[12] ),
    .C(\clkgen_inst.cnt_1s[19] ),
    .D(\clkgen_inst.cnt_1s[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_027_));
 sky130_fd_sc_hd__or4b_1 _135_ (.A(\clkgen_inst.cnt_1s[7] ),
    .B(_027_),
    .C(\clkgen_inst.cnt_1s[6] ),
    .D_N(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_028_));
 sky130_fd_sc_hd__or4_1 _136_ (.A(_020_),
    .B(_021_),
    .C(_024_),
    .D(_028_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_029_));
 sky130_fd_sc_hd__and2_1 _137_ (.A(net17),
    .B(_029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_030_));
 sky130_fd_sc_hd__nand2_1 _138_ (.A(\clkgen_inst.cnt_1s[6] ),
    .B(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_031_));
 sky130_fd_sc_hd__or2_1 _139_ (.A(\clkgen_inst.cnt_1s[6] ),
    .B(_019_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_032_));
 sky130_fd_sc_hd__and3_1 _140_ (.A(net10),
    .B(_031_),
    .C(_032_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[6] ));
 sky130_fd_sc_hd__and4_1 _141_ (.A(\clkgen_inst.cnt_1s[5] ),
    .B(\clkgen_inst.cnt_1s[4] ),
    .C(\clkgen_inst.cnt_1s[7] ),
    .D(\clkgen_inst.cnt_1s[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _142_ (.A(_016_),
    .B(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_034_));
 sky130_fd_sc_hd__a211oi_1 _143_ (.A1(_072_),
    .A2(_031_),
    .B1(_034_),
    .C1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n28_o[7] ));
 sky130_fd_sc_hd__and3_1 _144_ (.A(\clkgen_inst.cnt_1s[8] ),
    .B(_016_),
    .C(_033_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_035_));
 sky130_fd_sc_hd__o21ai_1 _145_ (.A1(net44),
    .A2(_034_),
    .B1(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _146_ (.A(_035_),
    .B(_036_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n28_o[8] ));
 sky130_fd_sc_hd__and2_1 _147_ (.A(\clkgen_inst.cnt_1s[9] ),
    .B(_035_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_037_));
 sky130_fd_sc_hd__o21ai_1 _148_ (.A1(\clkgen_inst.cnt_1s[9] ),
    .A2(_035_),
    .B1(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _149_ (.A(_037_),
    .B(_038_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n28_o[9] ));
 sky130_fd_sc_hd__o21ai_1 _150_ (.A1(\clkgen_inst.cnt_1s[10] ),
    .A2(_037_),
    .B1(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_039_));
 sky130_fd_sc_hd__a21oi_1 _151_ (.A1(net39),
    .A2(_037_),
    .B1(_039_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n28_o[10] ));
 sky130_fd_sc_hd__a31o_1 _152_ (.A1(\clkgen_inst.cnt_1s[9] ),
    .A2(\clkgen_inst.cnt_1s[10] ),
    .A3(_035_),
    .B1(\clkgen_inst.cnt_1s[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_040_));
 sky130_fd_sc_hd__and4_1 _153_ (.A(\clkgen_inst.cnt_1s[9] ),
    .B(\clkgen_inst.cnt_1s[8] ),
    .C(\clkgen_inst.cnt_1s[10] ),
    .D(\clkgen_inst.cnt_1s[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_041_));
 sky130_fd_sc_hd__and3_1 _154_ (.A(_016_),
    .B(_033_),
    .C(_041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_042_));
 sky130_fd_sc_hd__and3b_1 _155_ (.A_N(_042_),
    .B(net10),
    .C(_040_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[11] ));
 sky130_fd_sc_hd__and2_1 _156_ (.A(\clkgen_inst.cnt_1s[12] ),
    .B(_042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_043_));
 sky130_fd_sc_hd__or2_1 _157_ (.A(\clkgen_inst.cnt_1s[12] ),
    .B(_042_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_044_));
 sky130_fd_sc_hd__and3b_1 _158_ (.A_N(_043_),
    .B(_044_),
    .C(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[12] ));
 sky130_fd_sc_hd__and4_1 _159_ (.A(_016_),
    .B(_025_),
    .C(_033_),
    .D(_041_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_045_));
 sky130_fd_sc_hd__inv_2 _160_ (.A(_045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_046_));
 sky130_fd_sc_hd__o211a_1 _161_ (.A1(net42),
    .A2(_043_),
    .B1(_046_),
    .C1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[13] ));
 sky130_fd_sc_hd__or2_1 _162_ (.A(\clkgen_inst.cnt_1s[14] ),
    .B(_045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_047_));
 sky130_fd_sc_hd__o211a_1 _163_ (.A1(_073_),
    .A2(_046_),
    .B1(_047_),
    .C1(net10),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[14] ));
 sky130_fd_sc_hd__a21o_1 _164_ (.A1(\clkgen_inst.cnt_1s[14] ),
    .A2(_045_),
    .B1(\clkgen_inst.cnt_1s[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_048_));
 sky130_fd_sc_hd__and3_1 _165_ (.A(\clkgen_inst.cnt_1s[15] ),
    .B(\clkgen_inst.cnt_1s[14] ),
    .C(_045_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_049_));
 sky130_fd_sc_hd__and3b_1 _166_ (.A_N(_049_),
    .B(net18),
    .C(_048_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[15] ));
 sky130_fd_sc_hd__or2_1 _167_ (.A(\clkgen_inst.cnt_1s[16] ),
    .B(_049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_050_));
 sky130_fd_sc_hd__nand2_1 _168_ (.A(\clkgen_inst.cnt_1s[16] ),
    .B(_049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_051_));
 sky130_fd_sc_hd__and3_1 _169_ (.A(net10),
    .B(_050_),
    .C(_051_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[16] ));
 sky130_fd_sc_hd__a21oi_1 _170_ (.A1(\clkgen_inst.cnt_1s[16] ),
    .A2(_049_),
    .B1(\clkgen_inst.cnt_1s[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_052_));
 sky130_fd_sc_hd__a31o_1 _171_ (.A1(\clkgen_inst.cnt_1s[17] ),
    .A2(\clkgen_inst.cnt_1s[16] ),
    .A3(_049_),
    .B1(_071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_053_));
 sky130_fd_sc_hd__nor2_1 _172_ (.A(_052_),
    .B(_053_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n28_o[17] ));
 sky130_fd_sc_hd__a31o_1 _173_ (.A1(\clkgen_inst.cnt_1s[17] ),
    .A2(\clkgen_inst.cnt_1s[16] ),
    .A3(_049_),
    .B1(\clkgen_inst.cnt_1s[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_054_));
 sky130_fd_sc_hd__and4_1 _174_ (.A(\clkgen_inst.cnt_1s[17] ),
    .B(\clkgen_inst.cnt_1s[16] ),
    .C(\clkgen_inst.cnt_1s[18] ),
    .D(_049_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_055_));
 sky130_fd_sc_hd__and3b_1 _175_ (.A_N(_055_),
    .B(_030_),
    .C(_054_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[18] ));
 sky130_fd_sc_hd__and4_1 _176_ (.A(\clkgen_inst.cnt_1s[17] ),
    .B(\clkgen_inst.cnt_1s[16] ),
    .C(\clkgen_inst.cnt_1s[19] ),
    .D(\clkgen_inst.cnt_1s[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_056_));
 sky130_fd_sc_hd__and4_1 _177_ (.A(\clkgen_inst.cnt_1s[15] ),
    .B(\clkgen_inst.cnt_1s[14] ),
    .C(_045_),
    .D(_056_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_057_));
 sky130_fd_sc_hd__inv_2 _178_ (.A(_057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_058_));
 sky130_fd_sc_hd__o211a_1 _179_ (.A1(net43),
    .A2(_055_),
    .B1(_058_),
    .C1(_030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[19] ));
 sky130_fd_sc_hd__or2_1 _180_ (.A(\clkgen_inst.cnt_1s[20] ),
    .B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_059_));
 sky130_fd_sc_hd__nand2_1 _181_ (.A(\clkgen_inst.cnt_1s[20] ),
    .B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_060_));
 sky130_fd_sc_hd__and3_1 _182_ (.A(net10),
    .B(_059_),
    .C(_060_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[20] ));
 sky130_fd_sc_hd__a21o_1 _183_ (.A1(\clkgen_inst.cnt_1s[20] ),
    .A2(net11),
    .B1(\clkgen_inst.cnt_1s[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_061_));
 sky130_fd_sc_hd__nand2_1 _184_ (.A(_026_),
    .B(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_062_));
 sky130_fd_sc_hd__and3_1 _185_ (.A(net10),
    .B(_061_),
    .C(_062_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[21] ));
 sky130_fd_sc_hd__a21o_1 _186_ (.A1(_026_),
    .A2(net11),
    .B1(\clkgen_inst.cnt_1s[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_063_));
 sky130_fd_sc_hd__nand3_1 _187_ (.A(\clkgen_inst.cnt_1s[22] ),
    .B(_026_),
    .C(net11),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_064_));
 sky130_fd_sc_hd__and3_1 _188_ (.A(net10),
    .B(_063_),
    .C(_064_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[22] ));
 sky130_fd_sc_hd__and3_1 _189_ (.A(\clkgen_inst.cnt_1s[23] ),
    .B(\clkgen_inst.cnt_1s[22] ),
    .C(_026_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_065_));
 sky130_fd_sc_hd__a221oi_1 _190_ (.A1(_074_),
    .A2(_064_),
    .B1(_065_),
    .B2(net11),
    .C1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n28_o[23] ));
 sky130_fd_sc_hd__a21o_1 _191_ (.A1(net11),
    .A2(_065_),
    .B1(\clkgen_inst.cnt_1s[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_066_));
 sky130_fd_sc_hd__nand3_1 _192_ (.A(\clkgen_inst.cnt_1s[24] ),
    .B(net11),
    .C(_065_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_067_));
 sky130_fd_sc_hd__and3_1 _193_ (.A(net10),
    .B(_066_),
    .C(_067_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\clkgen_inst.n28_o[24] ));
 sky130_fd_sc_hd__a41o_1 _194_ (.A1(\clkgen_inst.cnt_1s[25] ),
    .A2(\clkgen_inst.cnt_1s[24] ),
    .A3(net11),
    .A4(_065_),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_068_));
 sky130_fd_sc_hd__a21oi_1 _195_ (.A1(_075_),
    .A2(_067_),
    .B1(_068_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\clkgen_inst.n28_o[25] ));
 sky130_fd_sc_hd__xor2_1 _196_ (.A(net40),
    .B(_029_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_069_));
 sky130_fd_sc_hd__nor2_1 _197_ (.A(net12),
    .B(_069_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_000_));
 sky130_fd_sc_hd__mux2_1 _198_ (.A0(htol_latched),
    .A1(net3),
    .S(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_001_));
 sky130_fd_sc_hd__a21oi_1 _199_ (.A1(_077_),
    .A2(_081_),
    .B1(net12),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(_070_));
 sky130_fd_sc_hd__o21a_1 _200_ (.A1(_077_),
    .A2(_081_),
    .B1(_070_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(_002_));
 sky130_fd_sc_hd__dfrtp_1 _201_ (.CLK(clknet_2_3__leaf_clk),
    .D(_000_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.htol_1s_toggle ));
 sky130_fd_sc_hd__dfrtp_2 _202_ (.CLK(clknet_2_3__leaf_clk),
    .D(_001_),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(htol_latched));
 sky130_fd_sc_hd__dfrtp_1 _203_ (.CLK(clknet_2_1__leaf_clk),
    .D(_002_),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.htol_1Mhz_toggle ));
 sky130_fd_sc_hd__dfrtp_1 _204_ (.CLK(clknet_2_1__leaf_clk),
    .D(\clkgen_inst.n30_o[0] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1m[0] ));
 sky130_fd_sc_hd__dfrtp_1 _205_ (.CLK(clknet_2_1__leaf_clk),
    .D(\clkgen_inst.n30_o[1] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1m[1] ));
 sky130_fd_sc_hd__dfrtp_1 _206_ (.CLK(clknet_2_0__leaf_clk),
    .D(\clkgen_inst.n30_o[2] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1m[2] ));
 sky130_fd_sc_hd__dfrtp_1 _207_ (.CLK(clknet_2_1__leaf_clk),
    .D(\clkgen_inst.n30_o[3] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1m[3] ));
 sky130_fd_sc_hd__dfrtp_1 _208_ (.CLK(clknet_2_1__leaf_clk),
    .D(\clkgen_inst.n30_o[4] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1m[4] ));
 sky130_fd_sc_hd__dfrtp_1 _209_ (.CLK(clknet_2_1__leaf_clk),
    .D(\clkgen_inst.n30_o[5] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1m[5] ));
 sky130_fd_sc_hd__dfrtp_2 _210_ (.CLK(clknet_2_3__leaf_clk),
    .D(\clkgen_inst.n28_o[0] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[0] ));
 sky130_fd_sc_hd__dfrtp_1 _211_ (.CLK(clknet_2_3__leaf_clk),
    .D(\clkgen_inst.n28_o[1] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[1] ));
 sky130_fd_sc_hd__dfrtp_1 _212_ (.CLK(clknet_2_3__leaf_clk),
    .D(\clkgen_inst.n28_o[2] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[2] ));
 sky130_fd_sc_hd__dfrtp_1 _213_ (.CLK(clknet_2_3__leaf_clk),
    .D(\clkgen_inst.n28_o[3] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[3] ));
 sky130_fd_sc_hd__dfrtp_1 _214_ (.CLK(clknet_2_3__leaf_clk),
    .D(\clkgen_inst.n28_o[4] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[4] ));
 sky130_fd_sc_hd__dfrtp_1 _215_ (.CLK(clknet_2_0__leaf_clk),
    .D(\clkgen_inst.n28_o[5] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[5] ));
 sky130_fd_sc_hd__dfrtp_1 _216_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[6] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[6] ));
 sky130_fd_sc_hd__dfrtp_1 _217_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[7] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[7] ));
 sky130_fd_sc_hd__dfrtp_1 _218_ (.CLK(clknet_2_3__leaf_clk),
    .D(\clkgen_inst.n28_o[8] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[8] ));
 sky130_fd_sc_hd__dfrtp_1 _219_ (.CLK(clknet_2_3__leaf_clk),
    .D(\clkgen_inst.n28_o[9] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[9] ));
 sky130_fd_sc_hd__dfrtp_1 _220_ (.CLK(clknet_2_3__leaf_clk),
    .D(\clkgen_inst.n28_o[10] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[10] ));
 sky130_fd_sc_hd__dfrtp_1 _221_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[11] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[11] ));
 sky130_fd_sc_hd__dfrtp_1 _222_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[12] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[12] ));
 sky130_fd_sc_hd__dfrtp_1 _223_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[13] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[13] ));
 sky130_fd_sc_hd__dfrtp_1 _224_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[14] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[14] ));
 sky130_fd_sc_hd__dfrtp_1 _225_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[15] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[15] ));
 sky130_fd_sc_hd__dfrtp_2 _226_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[16] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[16] ));
 sky130_fd_sc_hd__dfrtp_1 _227_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[17] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[17] ));
 sky130_fd_sc_hd__dfrtp_1 _228_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[18] ),
    .RESET_B(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[18] ));
 sky130_fd_sc_hd__dfrtp_1 _229_ (.CLK(clknet_2_2__leaf_clk),
    .D(\clkgen_inst.n28_o[19] ),
    .RESET_B(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[19] ));
 sky130_fd_sc_hd__dfrtp_1 _230_ (.CLK(clknet_2_0__leaf_clk),
    .D(\clkgen_inst.n28_o[20] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[20] ));
 sky130_fd_sc_hd__dfrtp_1 _231_ (.CLK(clknet_2_0__leaf_clk),
    .D(\clkgen_inst.n28_o[21] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[21] ));
 sky130_fd_sc_hd__dfrtp_1 _232_ (.CLK(clknet_2_0__leaf_clk),
    .D(\clkgen_inst.n28_o[22] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[22] ));
 sky130_fd_sc_hd__dfrtp_1 _233_ (.CLK(clknet_2_0__leaf_clk),
    .D(\clkgen_inst.n28_o[23] ),
    .RESET_B(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[23] ));
 sky130_fd_sc_hd__dfrtp_1 _234_ (.CLK(clknet_2_0__leaf_clk),
    .D(\clkgen_inst.n28_o[24] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[24] ));
 sky130_fd_sc_hd__dfrtp_1 _235_ (.CLK(clknet_2_0__leaf_clk),
    .D(\clkgen_inst.n28_o[25] ),
    .RESET_B(net13),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\clkgen_inst.cnt_1s[25] ));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net20));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net21));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net22));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net23));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net24));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net25));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net26));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net27));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net28));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net29));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net30));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net31));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net32));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net33));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net34));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net35));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net36));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_2 _254_ (.A(n55_o),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[0]));
 sky130_fd_sc_hd__buf_2 _255_ (.A(chain_out),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(uo_out[1]));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1000_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1000_inv_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1000_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1001_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1000_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1001_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1002_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1001_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1002_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1003_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1002_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1003_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1004_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1003_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1004_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1005_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1004_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1005_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1006_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1005_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1006_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1007_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1006_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1007_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1008_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1007_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1008_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1009_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1008_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1009_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n100_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n100_inv_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n100_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1010_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1009_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1010_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1011_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1010_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1011_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1012_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1011_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1012_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1013_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1012_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1013_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1014_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1013_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1014_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1015_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1014_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1015_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1016_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1015_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1016_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1017_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1016_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1017_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1018_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1017_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1018_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1019_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1018_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1019_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n101_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n100_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n101_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1020_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1019_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1020_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1021_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1020_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1021_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1022_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1021_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1022_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1023_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1022_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1023_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1024_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1023_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(chain_out));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n102_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n101_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n102_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n103_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n102_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n103_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n104_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n103_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n104_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n105_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n104_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n105_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n106_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n105_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n106_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n107_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n106_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n107_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n108_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n107_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n108_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n109_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n108_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n109_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n10_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n10_inv_inst.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n10_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n110_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n109_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n110_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n111_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n110_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n111_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n112_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n111_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n112_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n113_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n112_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n113_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n114_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n113_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n114_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n115_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n114_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n115_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n116_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n115_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n116_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n117_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n116_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n117_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n118_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n117_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n118_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n119_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n118_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n119_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n11_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n10_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n11_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n120_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n119_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n120_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n121_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n120_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n121_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n122_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n121_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n122_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n123_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n122_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n123_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n124_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n123_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n124_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n125_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n124_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n125_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n126_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n125_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n126_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n127_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n126_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n127_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n128_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n127_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n128_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n129_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n128_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n129_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n12_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n11_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n12_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n130_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n129_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n130_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n131_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n130_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n131_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n132_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n131_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n132_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n133_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n132_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n133_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n134_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n133_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n134_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n135_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n134_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n135_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n136_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n135_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n136_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n137_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n136_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n137_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n138_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n137_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n138_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n139_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n138_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n139_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n13_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n12_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n13_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n140_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n139_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n140_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n141_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n140_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n141_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n142_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n141_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n142_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n143_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n142_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n143_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n144_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n143_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n144_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n145_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n144_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n145_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n146_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n145_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n146_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n147_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n146_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n147_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n148_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n147_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n148_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n149_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n148_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n149_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n14_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n13_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n14_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n150_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n149_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n150_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n151_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n150_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n151_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n152_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n151_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n152_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n153_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n152_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n153_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n154_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n153_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n154_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n155_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n154_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n155_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n156_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n155_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n156_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n157_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n156_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n157_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n158_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n157_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n158_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n159_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n158_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n159_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n15_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n14_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n15_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n160_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n159_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n160_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n161_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n160_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n161_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n162_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n161_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n162_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n163_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n162_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n163_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n164_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n163_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n164_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n165_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n164_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n165_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n166_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n165_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n166_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n167_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n166_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n167_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n168_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n167_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n168_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n169_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n168_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n169_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n16_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n15_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n16_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n170_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n169_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n170_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n171_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n170_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n171_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n172_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n171_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n172_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n173_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n172_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n173_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n174_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n173_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n174_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n175_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n174_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n175_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n176_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n175_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n176_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n177_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n176_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n177_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n178_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n177_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n178_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n179_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n178_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n179_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n17_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n16_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n17_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n180_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n179_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n180_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n181_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n180_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n181_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n182_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n181_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n182_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n183_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n182_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n183_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n184_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n183_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n184_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n185_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n184_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n185_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n186_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n185_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n186_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n187_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n186_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n187_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n188_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n187_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n188_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n189_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n188_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n189_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n18_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n17_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n18_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n190_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n189_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n190_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n191_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n190_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n191_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n192_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n191_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n192_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n193_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n192_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n193_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n194_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n193_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n194_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n195_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n194_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n195_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n196_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n195_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n196_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n197_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n196_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n197_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n198_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n197_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n198_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n199_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n198_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n199_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n19_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n18_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n19_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n1_inv_inst.u_inv  (.A(net8),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n200_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n199_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n200_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n201_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n200_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n201_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n202_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n201_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n202_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n203_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n202_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n203_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n204_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n203_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n204_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n205_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n204_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n205_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n206_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n205_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n206_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n207_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n206_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n207_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n208_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n207_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n208_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n209_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n208_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n209_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n20_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n19_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n20_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n210_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n209_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n210_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n211_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n210_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n211_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n212_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n211_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n212_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n213_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n212_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n213_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n214_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n213_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n214_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n215_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n214_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n215_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n216_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n215_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n216_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n217_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n216_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n217_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n218_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n217_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n218_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n219_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n218_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n219_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n21_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n20_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n21_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n220_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n219_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n220_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n221_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n220_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n221_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n222_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n221_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n222_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n223_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n222_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n223_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n224_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n223_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n224_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n225_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n224_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n225_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n226_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n225_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n226_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n227_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n226_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n227_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n228_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n227_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n228_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n229_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n228_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n229_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n22_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n21_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n22_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n230_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n229_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n230_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n231_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n230_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n231_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n232_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n231_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n232_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n233_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n232_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n233_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n234_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n233_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n234_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n235_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n234_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n235_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n236_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n235_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n236_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n237_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n236_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n237_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n238_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n237_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n238_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n239_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n238_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n239_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n23_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n22_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n23_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n240_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n239_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n240_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n241_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n240_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n241_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n242_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n241_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n242_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n243_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n242_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n243_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n244_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n243_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n244_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n245_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n244_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n245_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n246_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n245_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n246_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n247_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n246_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n247_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n248_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n247_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n248_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n249_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n248_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n249_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n24_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n23_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n24_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n250_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n249_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n250_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n251_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n250_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n251_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n252_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n251_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n252_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n253_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n252_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n253_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n254_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n253_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n254_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n255_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n254_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n255_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n256_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n255_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n256_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n257_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n256_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n257_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n258_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n257_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n258_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n259_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n258_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n259_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n25_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n24_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n25_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n260_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n259_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n260_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n261_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n260_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n261_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n262_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n261_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n262_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n263_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n262_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n263_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n264_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n263_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n264_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n265_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n264_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n265_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n266_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n265_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n266_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n267_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n266_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n267_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n268_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n267_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n268_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n269_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n268_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n269_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n26_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n25_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n26_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n270_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n269_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n270_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n271_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n270_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n271_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n272_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n271_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n272_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n273_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n272_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n273_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n274_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n273_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n274_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n275_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n274_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n275_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n276_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n275_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n276_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n277_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n276_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n277_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n278_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n277_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n278_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n279_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n278_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n279_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n27_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n26_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n27_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n280_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n279_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n280_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n281_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n280_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n281_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n282_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n281_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n282_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n283_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n282_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n283_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n284_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n283_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n284_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n285_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n284_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n285_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n286_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n285_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n286_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n287_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n286_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n287_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n288_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n287_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n288_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n289_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n288_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n289_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n28_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n27_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n28_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n290_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n289_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n290_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n291_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n290_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n291_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n292_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n291_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n292_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n293_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n292_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n293_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n294_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n293_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n294_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n295_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n294_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n295_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n296_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n295_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n296_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n297_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n296_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n297_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n298_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n297_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n298_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n299_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n298_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n299_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n29_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n28_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n29_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n2_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n1_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n2_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n300_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n299_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n300_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n301_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n300_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n301_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n302_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n301_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n302_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n303_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n302_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n303_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n304_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n303_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n304_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n305_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n304_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n305_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n306_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n305_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n306_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n307_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n306_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n307_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n308_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n307_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n308_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n309_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n308_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n309_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n30_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n29_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n30_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n310_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n309_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n310_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n311_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n310_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n311_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n312_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n311_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n312_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n313_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n312_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n313_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n314_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n313_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n314_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n315_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n314_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n315_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n316_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n315_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n316_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n317_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n316_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n317_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n318_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n317_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n318_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n319_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n318_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n319_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n31_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n30_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n31_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n320_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n319_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n320_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n321_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n320_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n321_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n322_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n321_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n322_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n323_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n322_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n323_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n324_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n323_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n324_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n325_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n324_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n325_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n326_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n325_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n326_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n327_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n326_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n327_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n328_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n327_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n328_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n329_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n328_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n329_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n32_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n31_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n32_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n330_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n329_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n330_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n331_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n330_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n331_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n332_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n331_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n332_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n333_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n332_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n333_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n334_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n333_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n334_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n335_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n334_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n335_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n336_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n335_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n336_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n337_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n336_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n337_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n338_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n337_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n338_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n339_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n338_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n339_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n33_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n32_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n33_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n340_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n339_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n340_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n341_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n340_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n341_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n342_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n341_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n342_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n343_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n342_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n343_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n344_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n343_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n344_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n345_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n344_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n345_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n346_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n345_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n346_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n347_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n346_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n347_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n348_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n347_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n348_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n349_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n348_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n349_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n34_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n33_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n34_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n350_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n349_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n350_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n351_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n350_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n351_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n352_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n351_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n352_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n353_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n352_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n353_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n354_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n353_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n354_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n355_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n354_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n355_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n356_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n355_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n356_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n357_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n356_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n357_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n358_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n357_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n358_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n359_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n358_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n359_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n35_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n34_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n35_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n360_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n359_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n360_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n361_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n360_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n361_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n362_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n361_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n362_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n363_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n362_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n363_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n364_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n363_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n364_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n365_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n364_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n365_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n366_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n365_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n366_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n367_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n366_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n367_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n368_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n367_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n368_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n369_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n368_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n369_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n36_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n35_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n36_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n370_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n369_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n370_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n371_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n370_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n371_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n372_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n371_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n372_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n373_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n372_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n373_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n374_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n373_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n374_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n375_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n374_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n375_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n376_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n375_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n376_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n377_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n376_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n377_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n378_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n377_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n378_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n379_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n378_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n379_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n37_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n36_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n37_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n380_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n379_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n380_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n381_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n380_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n381_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n382_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n381_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n382_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n383_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n382_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n383_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n384_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n383_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n384_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n385_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n384_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n385_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n386_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n385_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n386_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n387_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n386_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n387_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n388_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n387_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n388_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n389_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n388_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n389_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n38_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n37_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n38_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n390_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n389_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n390_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n391_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n390_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n391_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n392_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n391_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n392_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n393_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n392_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n393_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n394_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n393_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n394_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n395_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n394_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n395_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n396_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n395_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n396_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n397_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n396_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n397_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n398_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n397_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n398_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n399_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n398_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n399_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n39_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n38_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n39_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n3_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n2_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n3_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n400_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n399_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n400_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n401_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n400_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n401_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n402_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n401_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n402_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n403_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n402_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n403_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n404_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n403_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n404_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n405_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n404_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n405_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n406_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n405_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n406_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n407_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n406_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n407_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n408_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n407_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n408_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n409_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n408_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n409_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n40_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n39_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n40_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n410_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n409_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n410_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n411_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n410_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n411_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n412_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n411_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n412_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n413_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n412_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n413_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n414_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n413_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n414_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n415_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n414_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n415_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n416_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n415_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n416_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n417_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n416_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n417_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n418_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n417_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n418_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n419_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n418_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n419_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n41_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n40_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n41_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n420_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n419_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n420_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n421_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n420_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n421_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n422_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n421_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n422_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n423_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n422_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n423_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n424_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n423_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n424_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n425_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n424_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n425_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n426_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n425_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n426_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n427_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n426_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n427_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n428_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n427_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n428_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n429_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n428_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n429_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n42_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n41_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n42_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n430_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n429_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n430_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n431_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n430_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n431_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n432_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n431_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n432_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n433_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n432_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n433_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n434_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n433_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n434_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n435_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n434_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n435_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n436_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n435_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n436_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n437_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n436_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n437_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n438_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n437_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n438_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n439_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n438_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n439_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n43_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n42_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n43_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n440_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n439_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n440_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n441_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n440_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n441_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n442_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n441_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n442_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n443_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n442_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n443_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n444_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n443_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n444_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n445_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n444_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n445_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n446_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n445_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n446_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n447_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n446_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n447_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n448_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n447_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n448_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n449_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n448_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n449_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n44_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n43_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n44_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n450_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n449_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n450_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n451_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n450_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n451_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n452_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n451_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n452_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n453_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n452_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n453_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n454_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n453_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n454_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n455_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n454_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n455_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n456_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n455_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n456_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n457_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n456_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n457_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n458_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n457_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n458_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n459_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n458_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n459_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n45_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n44_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n45_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n460_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n459_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n460_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n461_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n460_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n461_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n462_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n461_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n462_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n463_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n462_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n463_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n464_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n463_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n464_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n465_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n464_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n465_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n466_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n465_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n466_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n467_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n466_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n467_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n468_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n467_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n468_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n469_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n468_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n469_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n46_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n45_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n46_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n470_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n469_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n470_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n471_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n470_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n471_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n472_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n471_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n472_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n473_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n472_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n473_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n474_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n473_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n474_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n475_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n474_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n475_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n476_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n475_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n476_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n477_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n476_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n477_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n478_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n477_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n478_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n479_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n478_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n479_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n47_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n46_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n47_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n480_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n479_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n480_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n481_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n480_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n481_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n482_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n481_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n482_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n483_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n482_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n483_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n484_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n483_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n484_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n485_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n484_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n485_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n486_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n485_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n486_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n487_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n486_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n487_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n488_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n487_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n488_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n489_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n488_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n489_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n48_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n47_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n48_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n490_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n489_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n490_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n491_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n490_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n491_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n492_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n491_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n492_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n493_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n492_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n493_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n494_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n493_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n494_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n495_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n494_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n495_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n496_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n495_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n496_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n497_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n496_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n497_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n498_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n497_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n498_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n499_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n498_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n499_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n49_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n48_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n49_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n4_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n3_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n4_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n500_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n499_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n500_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n501_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n500_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n501_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n502_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n501_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n502_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n503_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n502_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n503_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n504_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n503_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n504_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n505_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n504_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n505_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n506_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n505_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n506_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n507_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n506_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n507_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n508_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n507_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n508_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n509_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n508_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n509_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n50_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n49_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n50_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n510_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n509_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n510_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n511_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n510_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n511_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n512_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n511_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.chain_mid ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n513_inv_inst.u_inv  (.A(\inverterchain_inst.chain_mid ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n513_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n514_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n513_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n514_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n515_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n514_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n515_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n516_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n515_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n516_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n517_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n516_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n517_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n518_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n517_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n518_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n519_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n518_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n519_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n51_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n50_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n51_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n520_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n519_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n520_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n521_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n520_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n521_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n522_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n521_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n522_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n523_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n522_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n523_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n524_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n523_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n524_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n525_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n524_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n525_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n526_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n525_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n526_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n527_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n526_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n527_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n528_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n527_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n528_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n529_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n528_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n529_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n52_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n51_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n52_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n530_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n529_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n530_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n531_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n530_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n531_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n532_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n531_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n532_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n533_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n532_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n533_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n534_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n533_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n534_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n535_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n534_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n535_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n536_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n535_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n536_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n537_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n536_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n537_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n538_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n537_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n538_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n539_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n538_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n539_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n53_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n52_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n53_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n540_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n539_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n540_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n541_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n540_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n541_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n542_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n541_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n542_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n543_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n542_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n543_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n544_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n543_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n544_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n545_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n544_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n545_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n546_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n545_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n546_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n547_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n546_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n547_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n548_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n547_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n548_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n549_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n548_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n549_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n54_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n53_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n54_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n550_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n549_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n550_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n551_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n550_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n551_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n552_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n551_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n552_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n553_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n552_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n553_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n554_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n553_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n554_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n555_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n554_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n555_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n556_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n555_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n556_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n557_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n556_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n557_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n558_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n557_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n558_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n559_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n558_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n559_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n55_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n54_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n55_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n560_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n559_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n560_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n561_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n560_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n561_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n562_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n561_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n562_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n563_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n562_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n563_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n564_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n563_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n564_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n565_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n564_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n565_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n566_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n565_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n566_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n567_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n566_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n567_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n568_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n567_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n568_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n569_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n568_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n569_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n56_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n55_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n56_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n570_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n569_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n570_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n571_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n570_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n571_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n572_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n571_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n572_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n573_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n572_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n573_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n574_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n573_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n574_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n575_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n574_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n575_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n576_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n575_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n576_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n577_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n576_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n577_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n578_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n577_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n578_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n579_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n578_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n579_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n57_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n56_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n57_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n580_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n579_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n580_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n581_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n580_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n581_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n582_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n581_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n582_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n583_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n582_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n583_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n584_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n583_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n584_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n585_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n584_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n585_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n586_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n585_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n586_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n587_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n586_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n587_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n588_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n587_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n588_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n589_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n588_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n589_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n58_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n57_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n58_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n590_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n589_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n590_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n591_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n590_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n591_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n592_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n591_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n592_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n593_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n592_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n593_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n594_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n593_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n594_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n595_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n594_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n595_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n596_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n595_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n596_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n597_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n596_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n597_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n598_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n597_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n598_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n599_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n598_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n599_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n59_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n58_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n59_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n5_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n4_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n5_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n600_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n599_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n600_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n601_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n600_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n601_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n602_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n601_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n602_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n603_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n602_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n603_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n604_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n603_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n604_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n605_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n604_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n605_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n606_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n605_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n606_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n607_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n606_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n607_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n608_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n607_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n608_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n609_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n608_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n609_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n60_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n59_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n60_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n610_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n609_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n610_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n611_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n610_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n611_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n612_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n611_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n612_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n613_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n612_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n613_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n614_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n613_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n614_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n615_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n614_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n615_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n616_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n615_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n616_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n617_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n616_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n617_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n618_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n617_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n618_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n619_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n618_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n619_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n61_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n60_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n61_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n620_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n619_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n620_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n621_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n620_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n621_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n622_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n621_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n622_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n623_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n622_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n623_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n624_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n623_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n624_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n625_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n624_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n625_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n626_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n625_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n626_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n627_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n626_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n627_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n628_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n627_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n628_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n629_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n628_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n629_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n62_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n61_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n62_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n630_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n629_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n630_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n631_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n630_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n631_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n632_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n631_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n632_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n633_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n632_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n633_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n634_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n633_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n634_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n635_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n634_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n635_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n636_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n635_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n636_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n637_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n636_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n637_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n638_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n637_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n638_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n639_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n638_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n639_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n63_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n62_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n63_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n640_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n639_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n640_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n641_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n640_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n641_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n642_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n641_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n642_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n643_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n642_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n643_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n644_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n643_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n644_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n645_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n644_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n645_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n646_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n645_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n646_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n647_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n646_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n647_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n648_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n647_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n648_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n649_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n648_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n649_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n64_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n63_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n64_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n650_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n649_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n650_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n651_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n650_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n651_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n652_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n651_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n652_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n653_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n652_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n653_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n654_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n653_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n654_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n655_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n654_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n655_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n656_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n655_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n656_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n657_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n656_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n657_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n658_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n657_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n658_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n659_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n658_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n659_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n65_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n64_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n65_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n660_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n659_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n660_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n661_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n660_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n661_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n662_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n661_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n662_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n663_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n662_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n663_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n664_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n663_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n664_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n665_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n664_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n665_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n666_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n665_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n666_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n667_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n666_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n667_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n668_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n667_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n668_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n669_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n668_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n669_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n66_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n65_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n66_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n670_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n669_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n670_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n671_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n670_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n671_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n672_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n671_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n672_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n673_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n672_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n673_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n674_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n673_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n674_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n675_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n674_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n675_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n676_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n675_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n676_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n677_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n676_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n677_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n678_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n677_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n678_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n679_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n678_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n679_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n67_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n66_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n67_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n680_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n679_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n680_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n681_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n680_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n681_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n682_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n681_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n682_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n683_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n682_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n683_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n684_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n683_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n684_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n685_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n684_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n685_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n686_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n685_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n686_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n687_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n686_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n687_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n688_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n687_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n688_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n689_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n688_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n689_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n68_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n67_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n68_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n690_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n689_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n690_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n691_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n690_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n691_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n692_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n691_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n692_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n693_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n692_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n693_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n694_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n693_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n694_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n695_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n694_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n695_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n696_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n695_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n696_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n697_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n696_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n697_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n698_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n697_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n698_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n699_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n698_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n699_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n69_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n68_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n69_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n6_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n5_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n6_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n700_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n699_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n700_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n701_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n700_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n701_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n702_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n701_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n702_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n703_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n702_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n703_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n704_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n703_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n704_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n705_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n704_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n705_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n706_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n705_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n706_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n707_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n706_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n707_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n708_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n707_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n708_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n709_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n708_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n709_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n70_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n69_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n70_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n710_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n709_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n710_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n711_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n710_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n711_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n712_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n711_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n712_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n713_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n712_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n713_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n714_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n713_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n714_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n715_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n714_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n715_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n716_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n715_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n716_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n717_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n716_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n717_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n718_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n717_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n718_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n719_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n718_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n719_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n71_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n70_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n71_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n720_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n719_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n720_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n721_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n720_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n721_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n722_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n721_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n722_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n723_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n722_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n723_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n724_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n723_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n724_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n725_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n724_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n725_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n726_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n725_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n726_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n727_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n726_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n727_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n728_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n727_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n728_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n729_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n728_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n729_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n72_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n71_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n72_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n730_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n729_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n730_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n731_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n730_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n731_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n732_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n731_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n732_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n733_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n732_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n733_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n734_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n733_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n734_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n735_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n734_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n735_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n736_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n735_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n736_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n737_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n736_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n737_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n738_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n737_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n738_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n739_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n738_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n739_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n73_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n72_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n73_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n740_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n739_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n740_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n741_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n740_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n741_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n742_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n741_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n742_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n743_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n742_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n743_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n744_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n743_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n744_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n745_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n744_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n745_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n746_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n745_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n746_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n747_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n746_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n747_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n748_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n747_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n748_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n749_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n748_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n749_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n74_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n73_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n74_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n750_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n749_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n750_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n751_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n750_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n751_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n752_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n751_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n752_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n753_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n752_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n753_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n754_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n753_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n754_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n755_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n754_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n755_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n756_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n755_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n756_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n757_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n756_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n757_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n758_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n757_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n758_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n759_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n758_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n759_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n75_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n74_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n75_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n760_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n759_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n760_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n761_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n760_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n761_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n762_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n761_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n762_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n763_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n762_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n763_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n764_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n763_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n764_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n765_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n764_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n765_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n766_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n765_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n766_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n767_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n766_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n767_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n768_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n767_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.chain_3q ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n769_inv_inst.u_inv  (.A(\inverterchain_inst.chain_3q ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n769_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n76_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n75_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n76_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n770_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n769_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n770_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n771_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n770_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n771_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n772_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n771_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n772_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n773_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n772_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n773_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n774_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n773_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n774_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n775_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n774_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n775_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n776_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n775_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n776_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n777_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n776_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n777_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n778_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n777_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n778_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n779_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n778_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n779_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n77_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n76_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n77_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n780_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n779_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n780_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n781_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n780_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n781_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n782_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n781_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n782_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n783_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n782_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n783_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n784_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n783_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n784_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n785_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n784_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n785_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n786_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n785_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n786_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n787_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n786_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n787_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n788_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n787_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n788_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n789_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n788_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n789_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n78_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n77_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n78_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n790_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n789_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n790_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n791_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n790_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n791_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n792_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n791_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n792_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n793_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n792_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n793_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n794_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n793_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n794_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n795_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n794_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n795_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n796_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n795_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n796_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n797_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n796_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n797_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n798_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n797_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n798_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n799_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n798_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n799_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n79_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n78_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n79_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n7_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n6_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n7_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n800_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n799_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n800_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n801_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n800_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n801_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n802_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n801_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n802_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n803_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n802_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n803_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n804_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n803_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n804_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n805_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n804_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n805_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n806_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n805_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n806_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n807_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n806_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n807_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n808_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n807_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n808_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n809_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n808_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n809_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n80_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n79_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n80_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n810_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n809_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n810_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n811_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n810_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n811_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n812_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n811_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n812_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n813_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n812_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n813_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n814_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n813_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n814_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n815_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n814_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n815_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n816_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n815_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n816_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n817_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n816_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n817_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n818_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n817_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n818_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n819_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n818_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n819_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n81_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n80_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n81_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n820_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n819_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n820_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n821_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n820_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n821_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n822_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n821_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n822_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n823_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n822_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n823_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n824_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n823_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n824_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n825_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n824_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n825_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n826_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n825_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n826_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n827_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n826_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n827_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n828_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n827_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n828_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n829_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n828_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n829_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n82_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n81_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n82_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n830_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n829_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n830_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n831_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n830_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n831_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n832_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n831_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n832_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n833_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n832_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n833_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n834_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n833_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n834_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n835_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n834_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n835_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n836_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n835_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n836_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n837_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n836_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n837_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n838_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n837_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n838_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n839_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n838_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n839_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n83_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n82_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n83_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n840_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n839_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n840_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n841_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n840_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n841_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n842_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n841_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n842_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n843_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n842_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n843_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n844_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n843_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n844_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n845_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n844_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n845_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n846_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n845_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n846_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n847_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n846_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n847_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n848_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n847_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n848_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n849_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n848_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n849_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n84_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n83_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n84_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n850_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n849_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n850_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n851_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n850_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n851_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n852_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n851_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n852_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n853_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n852_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n853_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n854_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n853_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n854_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n855_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n854_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n855_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n856_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n855_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n856_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n857_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n856_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n857_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n858_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n857_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n858_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n859_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n858_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n859_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n85_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n84_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n85_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n860_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n859_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n860_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n861_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n860_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n861_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n862_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n861_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n862_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n863_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n862_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n863_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n864_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n863_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n864_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n865_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n864_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n865_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n866_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n865_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n866_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n867_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n866_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n867_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n868_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n867_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n868_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n869_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n868_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n869_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n86_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n85_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n86_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n870_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n869_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n870_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n871_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n870_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n871_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n872_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n871_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n872_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n873_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n872_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n873_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n874_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n873_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n874_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n875_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n874_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n875_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n876_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n875_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n876_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n877_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n876_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n877_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n878_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n877_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n878_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n879_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n878_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n879_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n87_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n86_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n87_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n880_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n879_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n880_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n881_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n880_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n881_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n882_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n881_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n882_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n883_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n882_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n883_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n884_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n883_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n884_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n885_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n884_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n885_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n886_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n885_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n886_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n887_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n886_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n887_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n888_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n887_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n888_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n889_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n888_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n889_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n88_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n87_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n88_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n890_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n889_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n890_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n891_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n890_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n891_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n892_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n891_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n892_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n893_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n892_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n893_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n894_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n893_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n894_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n895_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n894_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n895_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n896_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n895_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n896_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n897_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n896_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n897_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n898_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n897_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n898_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n899_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n898_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n899_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n89_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n88_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n89_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n8_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n7_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n8_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n900_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n899_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n900_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n901_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n900_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n901_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n902_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n901_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n902_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n903_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n902_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n903_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n904_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n903_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n904_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n905_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n904_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n905_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n906_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n905_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n906_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n907_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n906_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n907_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n908_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n907_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n908_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n909_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n908_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n909_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n90_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n89_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n90_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n910_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n909_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n910_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n911_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n910_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n911_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n912_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n911_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n912_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n913_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n912_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n913_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n914_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n913_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n914_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n915_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n914_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n915_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n916_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n915_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n916_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n917_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n916_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n917_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n918_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n917_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n918_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n919_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n918_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n919_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n91_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n90_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n91_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n920_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n919_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n920_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n921_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n920_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n921_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n922_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n921_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n922_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n923_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n922_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n923_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n924_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n923_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n924_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n925_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n924_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n925_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n926_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n925_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n926_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n927_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n926_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n927_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n928_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n927_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n928_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n929_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n928_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n929_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n92_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n91_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n92_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n930_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n929_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n930_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n931_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n930_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n931_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n932_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n931_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n932_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n933_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n932_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n933_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n934_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n933_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n934_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n935_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n934_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n935_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n936_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n935_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n936_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n937_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n936_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n937_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n938_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n937_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n938_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n939_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n938_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n939_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n93_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n92_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n93_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n940_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n939_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n940_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n941_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n940_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n941_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n942_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n941_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n942_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n943_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n942_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n943_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n944_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n943_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n944_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n945_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n944_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n945_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n946_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n945_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n946_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n947_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n946_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n947_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n948_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n947_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n948_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n949_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n948_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n949_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n94_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n93_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n94_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n950_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n949_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n950_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n951_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n950_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n951_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n952_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n951_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n952_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n953_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n952_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n953_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n954_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n953_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n954_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n955_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n954_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n955_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n956_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n955_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n956_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n957_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n956_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n957_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n958_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n957_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n958_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n959_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n958_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n959_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n95_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n94_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n95_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n960_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n959_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n960_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n961_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n960_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n961_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n962_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n961_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n962_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n963_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n962_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n963_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n964_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n963_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n964_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n965_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n964_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n965_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n966_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n965_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n966_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n967_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n966_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n967_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n968_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n967_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n968_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n969_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n968_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n969_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n96_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n95_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n96_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n970_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n969_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n970_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n971_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n970_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n971_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n972_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n971_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n972_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n973_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n972_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n973_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n974_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n973_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n974_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n975_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n974_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n975_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n976_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n975_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n976_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n977_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n976_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n977_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n978_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n977_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n978_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n979_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n978_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n979_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n97_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n96_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n97_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n980_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n979_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n980_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n981_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n980_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n981_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n982_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n981_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n982_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n983_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n982_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n983_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n984_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n983_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n984_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n985_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n984_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n985_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n986_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n985_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n986_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n987_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n986_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n987_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n988_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n987_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n988_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n989_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n988_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n989_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n98_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n97_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n98_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n990_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n989_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n990_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n991_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n990_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n991_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n992_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n991_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n992_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n993_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n992_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n993_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n994_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n993_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n994_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n995_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n994_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n995_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n996_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n995_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n996_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n997_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n996_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n997_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n998_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n997_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n998_inv_inst.Y ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n999_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n998_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n1000_inv_inst.A ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n99_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n98_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n100_inv_inst.A ));
 sky130_fd_sc_hd__inv_1 \inverterchain_inst.gen_inv_n9_inv_inst.u_inv  (.A(\inverterchain_inst.gen_inv_n8_inv_inst.Y ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\inverterchain_inst.gen_inv_n10_inv_inst.A ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ena),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(rst_n),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(uio_in[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(uio_in[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(uio_in[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(uio_in[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(uio_in[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(uio_in[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(uio_in[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 fanout10 (.A(_030_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__buf_2 fanout11 (.A(_057_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(_071_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 fanout14 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(net2),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 fanout18 (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__conb_1 tt_um_technology_characterization_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net19));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_2_0__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__bufinv_16 clkload1 (.A(clknet_2_1__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload2 (.A(clknet_2_3__leaf_clk),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\clkgen_inst.cnt_1m[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\clkgen_inst.cnt_1s[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\clkgen_inst.cnt_1s[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\clkgen_inst.htol_1s_toggle ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\clkgen_inst.cnt_1m[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\clkgen_inst.cnt_1s[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\clkgen_inst.cnt_1s[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\clkgen_inst.cnt_1s[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\clkgen_inst.cnt_1s[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\clkgen_inst.cnt_1s[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\clkgen_inst.cnt_1s[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\clkgen_inst.cnt_1m[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\clkgen_inst.cnt_1s[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_148 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_1_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_131 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_155 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_1_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_1_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_157 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_2_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_3_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_3_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_3_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_4_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_4_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_4_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_147 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_5_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_184 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_196 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_5_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_234 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_246 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_258 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_5_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_162 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_174 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_6_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_6_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_7_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_7_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_7_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_133 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_7_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_7_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_251 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_8_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_157 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_8_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_215 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_8_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_9_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_9_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_151 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_9_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_9_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_9_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_250 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_262 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_10_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_10_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_217 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_10_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_10_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_10_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_11_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_88 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_100 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_152 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_11_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_11_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_251 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_11_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_11_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_12_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_114 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_126 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_12_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_12_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_12_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_12_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_12_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_12_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_13_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_13_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_13_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_143 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_13_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_13_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_14_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_114 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_14_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_158 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_170 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_14_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_14_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_271 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_283 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_14_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_318 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_14_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_15_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_75 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_15_87 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_15_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_154 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_15_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_15_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_15_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_287 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_15_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_315 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_15_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_16_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_16_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_16_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_229 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_16_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_312 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_16_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_17_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_60 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_72 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_17_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_17_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_142 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_154 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_17_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_202 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_17_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_228 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_17_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_303 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_315 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_17_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_18_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_18_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_227 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_18_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_18_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_19_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_19_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_19_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_19_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_284 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_19_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_314 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_19_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_20_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_20_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_20_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_259 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_280 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_323 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_21_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_21_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_21_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_138 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_21_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_192 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_204 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_21_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_21_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_21_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_22_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_22_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_63 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_22_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_106 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_22_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_179 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_22_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_207 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_22_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_234 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_22_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_23_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_127 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_23_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_301 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_316 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_23_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_51 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_63 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_24_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_24_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_106 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_118 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_24_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_151 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_163 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_24_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_206 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_24_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_238 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_24_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_24_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_24_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_24_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_25_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_25_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_25_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_264 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_25_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_26_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_67 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_26_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_151 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_26_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_217 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_26_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_239 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_26_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_322 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_26_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_27_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_62 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_27_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_120 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_132 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_27_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_240 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_27_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_28_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_88 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_28_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_279 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_28_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_28_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_29_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_63 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_29_75 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_29_87 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_29_99 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_29_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_135 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_29_147 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_29_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_30_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_30_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_47 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_30_59 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_30_71 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_30_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_30_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_30_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_30_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_316 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_30_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_67 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_79 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_31_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_31_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_135 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_31_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_31_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_31_285 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_31_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_32_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_49 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_32_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_32_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_32_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_33_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_33_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_71 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_33_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_33_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_323 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_34_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_34_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_34_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_34_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_34_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_35_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_35_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_35_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_35_301 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_35_313 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_35_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_36_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_36_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_36_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_36_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_36_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_238 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_36_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_280 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_292 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_36_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_36_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_37_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_63 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_75 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_87 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_99 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_37_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_37_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_37_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_38_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_38_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_38_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_38_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_38_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_316 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_38_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 assign uio_oe[0] = net19;
 assign uio_oe[1] = net20;
 assign uio_oe[2] = net21;
 assign uio_oe[3] = net22;
 assign uio_oe[4] = net23;
 assign uio_oe[5] = net24;
 assign uio_oe[6] = net25;
 assign uio_oe[7] = net26;
 assign uio_out[0] = net27;
 assign uio_out[1] = net28;
 assign uio_out[2] = net29;
 assign uio_out[3] = net30;
 assign uio_out[4] = net31;
 assign uio_out[5] = net32;
 assign uio_out[6] = net33;
 assign uio_out[7] = net34;
 assign uo_out[2] = net35;
 assign uo_out[3] = net36;
endmodule
